--Connor Murphy
--Section 11092

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity shift_left_2 is
    port (
        input : in std_logic_vector(31 downto 0);
        output : out std_logic_vector(31 downto 0)
    );
end shift_left_2;

architecture behavioral of shift_left_2 is
    -- Placeholder
begin
    -- Placeholder
end behavioral;