--Connor Murphy
--Section 11092

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity shift_left_2_28bit is
    port (
        input : in std_logic_vector(25 downto 0);
        output : out std_logic_vector(27 downto 0)
    );
end shift_left_2_28bit;

architecture behavioral of shift_left_2_28bit is
    -- Placeholder
begin
    -- Placeholder
end behavioral;